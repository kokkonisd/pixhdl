library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity W150_Adder is
Port (  CLK, RST, WE : in STD_LOGIC;
        Bias     : in STD_LOGIC_VECTOR (31 downto 0);
        Float001 : in STD_LOGIC_VECTOR (31 downto 0);
        Float002 : in STD_LOGIC_VECTOR (31 downto 0);
        Float003 : in STD_LOGIC_VECTOR (31 downto 0);
        Float004 : in STD_LOGIC_VECTOR (31 downto 0);
        Float005 : in STD_LOGIC_VECTOR (31 downto 0);
        Float006 : in STD_LOGIC_VECTOR (31 downto 0);
        Float007 : in STD_LOGIC_VECTOR (31 downto 0);
        Float008 : in STD_LOGIC_VECTOR (31 downto 0);
        Float009 : in STD_LOGIC_VECTOR (31 downto 0);
        Float010 : in STD_LOGIC_VECTOR (31 downto 0);
        Float011 : in STD_LOGIC_VECTOR (31 downto 0);
        Float012 : in STD_LOGIC_VECTOR (31 downto 0);
        Float013 : in STD_LOGIC_VECTOR (31 downto 0);
        Float014 : in STD_LOGIC_VECTOR (31 downto 0);
        Float015 : in STD_LOGIC_VECTOR (31 downto 0);
        Float016 : in STD_LOGIC_VECTOR (31 downto 0);
        Float017 : in STD_LOGIC_VECTOR (31 downto 0);
        Float018 : in STD_LOGIC_VECTOR (31 downto 0);
        Float019 : in STD_LOGIC_VECTOR (31 downto 0);
        Float020 : in STD_LOGIC_VECTOR (31 downto 0);
        Float021 : in STD_LOGIC_VECTOR (31 downto 0);
        Float022 : in STD_LOGIC_VECTOR (31 downto 0);
        Float023 : in STD_LOGIC_VECTOR (31 downto 0);
        Float024 : in STD_LOGIC_VECTOR (31 downto 0);
        Float025 : in STD_LOGIC_VECTOR (31 downto 0);
        Float026 : in STD_LOGIC_VECTOR (31 downto 0);
        Float027 : in STD_LOGIC_VECTOR (31 downto 0);
        Float028 : in STD_LOGIC_VECTOR (31 downto 0);
        Float029 : in STD_LOGIC_VECTOR (31 downto 0);
        Float030 : in STD_LOGIC_VECTOR (31 downto 0);
        Float031 : in STD_LOGIC_VECTOR (31 downto 0);
        Float032 : in STD_LOGIC_VECTOR (31 downto 0);
        Float033 : in STD_LOGIC_VECTOR (31 downto 0);
        Float034 : in STD_LOGIC_VECTOR (31 downto 0);
        Float035 : in STD_LOGIC_VECTOR (31 downto 0);
        Float036 : in STD_LOGIC_VECTOR (31 downto 0);
        Float037 : in STD_LOGIC_VECTOR (31 downto 0);
        Float038 : in STD_LOGIC_VECTOR (31 downto 0);
        Float039 : in STD_LOGIC_VECTOR (31 downto 0);
        Float040 : in STD_LOGIC_VECTOR (31 downto 0);
        Float041 : in STD_LOGIC_VECTOR (31 downto 0);
        Float042 : in STD_LOGIC_VECTOR (31 downto 0);
        Float043 : in STD_LOGIC_VECTOR (31 downto 0);
        Float044 : in STD_LOGIC_VECTOR (31 downto 0);
        Float045 : in STD_LOGIC_VECTOR (31 downto 0);
        Float046 : in STD_LOGIC_VECTOR (31 downto 0);
        Float047 : in STD_LOGIC_VECTOR (31 downto 0);
        Float048 : in STD_LOGIC_VECTOR (31 downto 0);
        Float049 : in STD_LOGIC_VECTOR (31 downto 0);
        Float050 : in STD_LOGIC_VECTOR (31 downto 0);
        Float051 : in STD_LOGIC_VECTOR (31 downto 0);
        Float052 : in STD_LOGIC_VECTOR (31 downto 0);
        Float053 : in STD_LOGIC_VECTOR (31 downto 0);
        Float054 : in STD_LOGIC_VECTOR (31 downto 0);
        Float055 : in STD_LOGIC_VECTOR (31 downto 0);
        Float056 : in STD_LOGIC_VECTOR (31 downto 0);
        Float057 : in STD_LOGIC_VECTOR (31 downto 0);
        Float058 : in STD_LOGIC_VECTOR (31 downto 0);
        Float059 : in STD_LOGIC_VECTOR (31 downto 0);
        Float060 : in STD_LOGIC_VECTOR (31 downto 0);
        Float061 : in STD_LOGIC_VECTOR (31 downto 0);
        Float062 : in STD_LOGIC_VECTOR (31 downto 0);
        Float063 : in STD_LOGIC_VECTOR (31 downto 0);
        Float064 : in STD_LOGIC_VECTOR (31 downto 0);
        Float065 : in STD_LOGIC_VECTOR (31 downto 0);
        Float066 : in STD_LOGIC_VECTOR (31 downto 0);
        Float067 : in STD_LOGIC_VECTOR (31 downto 0);
        Float068 : in STD_LOGIC_VECTOR (31 downto 0);
        Float069 : in STD_LOGIC_VECTOR (31 downto 0);
        Float070 : in STD_LOGIC_VECTOR (31 downto 0);
        Float071 : in STD_LOGIC_VECTOR (31 downto 0);
        Float072 : in STD_LOGIC_VECTOR (31 downto 0);
        Float073 : in STD_LOGIC_VECTOR (31 downto 0);
        Float074 : in STD_LOGIC_VECTOR (31 downto 0);
        Float075 : in STD_LOGIC_VECTOR (31 downto 0);
        Float076 : in STD_LOGIC_VECTOR (31 downto 0);
        Float077 : in STD_LOGIC_VECTOR (31 downto 0);
        Float078 : in STD_LOGIC_VECTOR (31 downto 0);
        Float079 : in STD_LOGIC_VECTOR (31 downto 0);
        Float080 : in STD_LOGIC_VECTOR (31 downto 0);
        Float081 : in STD_LOGIC_VECTOR (31 downto 0);
        Float082 : in STD_LOGIC_VECTOR (31 downto 0);
        Float083 : in STD_LOGIC_VECTOR (31 downto 0);
        Float084 : in STD_LOGIC_VECTOR (31 downto 0);
        Float085 : in STD_LOGIC_VECTOR (31 downto 0);
        Float086 : in STD_LOGIC_VECTOR (31 downto 0);
        Float087 : in STD_LOGIC_VECTOR (31 downto 0);
        Float088 : in STD_LOGIC_VECTOR (31 downto 0);
        Float089 : in STD_LOGIC_VECTOR (31 downto 0);
        Float090 : in STD_LOGIC_VECTOR (31 downto 0);
        Float091 : in STD_LOGIC_VECTOR (31 downto 0);
        Float092 : in STD_LOGIC_VECTOR (31 downto 0);
        Float093 : in STD_LOGIC_VECTOR (31 downto 0);
        Float094 : in STD_LOGIC_VECTOR (31 downto 0);
        Float095 : in STD_LOGIC_VECTOR (31 downto 0);
        Float096 : in STD_LOGIC_VECTOR (31 downto 0);
        Float097 : in STD_LOGIC_VECTOR (31 downto 0);
        Float098 : in STD_LOGIC_VECTOR (31 downto 0);
        Float099 : in STD_LOGIC_VECTOR (31 downto 0);
        Float100 : in STD_LOGIC_VECTOR (31 downto 0);
        Float101 : in STD_LOGIC_VECTOR (31 downto 0);
        Float102 : in STD_LOGIC_VECTOR (31 downto 0);
        Float103 : in STD_LOGIC_VECTOR (31 downto 0);
        Float104 : in STD_LOGIC_VECTOR (31 downto 0);
        Float105 : in STD_LOGIC_VECTOR (31 downto 0);
        Float106 : in STD_LOGIC_VECTOR (31 downto 0);
        Float107 : in STD_LOGIC_VECTOR (31 downto 0);
        Float108 : in STD_LOGIC_VECTOR (31 downto 0);
        Float109 : in STD_LOGIC_VECTOR (31 downto 0);
        Float110 : in STD_LOGIC_VECTOR (31 downto 0);
        Float111 : in STD_LOGIC_VECTOR (31 downto 0);
        Float112 : in STD_LOGIC_VECTOR (31 downto 0);
        Float113 : in STD_LOGIC_VECTOR (31 downto 0);
        Float114 : in STD_LOGIC_VECTOR (31 downto 0);
        Float115 : in STD_LOGIC_VECTOR (31 downto 0);
        Float116 : in STD_LOGIC_VECTOR (31 downto 0);
        Float117 : in STD_LOGIC_VECTOR (31 downto 0);
        Float118 : in STD_LOGIC_VECTOR (31 downto 0);
        Float119 : in STD_LOGIC_VECTOR (31 downto 0);
        Float120 : in STD_LOGIC_VECTOR (31 downto 0);
        Float121 : in STD_LOGIC_VECTOR (31 downto 0);
        Float122 : in STD_LOGIC_VECTOR (31 downto 0);
        Float123 : in STD_LOGIC_VECTOR (31 downto 0);
        Float124 : in STD_LOGIC_VECTOR (31 downto 0);
        Float125 : in STD_LOGIC_VECTOR (31 downto 0);
        Float126 : in STD_LOGIC_VECTOR (31 downto 0);
        Float127 : in STD_LOGIC_VECTOR (31 downto 0);
        Float128 : in STD_LOGIC_VECTOR (31 downto 0);
        Float129 : in STD_LOGIC_VECTOR (31 downto 0);
        Float130 : in STD_LOGIC_VECTOR (31 downto 0);
        Float131 : in STD_LOGIC_VECTOR (31 downto 0);
        Float132 : in STD_LOGIC_VECTOR (31 downto 0);
        Float133 : in STD_LOGIC_VECTOR (31 downto 0);
        Float134 : in STD_LOGIC_VECTOR (31 downto 0);
        Float135 : in STD_LOGIC_VECTOR (31 downto 0);
        Float136 : in STD_LOGIC_VECTOR (31 downto 0);
        Float137 : in STD_LOGIC_VECTOR (31 downto 0);
        Float138 : in STD_LOGIC_VECTOR (31 downto 0);
        Float139 : in STD_LOGIC_VECTOR (31 downto 0);
        Float140 : in STD_LOGIC_VECTOR (31 downto 0);
        Float141 : in STD_LOGIC_VECTOR (31 downto 0);
        Float142 : in STD_LOGIC_VECTOR (31 downto 0);
        Float143 : in STD_LOGIC_VECTOR (31 downto 0);
        Float144 : in STD_LOGIC_VECTOR (31 downto 0);
        Float145 : in STD_LOGIC_VECTOR (31 downto 0);
        Float146 : in STD_LOGIC_VECTOR (31 downto 0);
        Float147 : in STD_LOGIC_VECTOR (31 downto 0);
        Float148 : in STD_LOGIC_VECTOR (31 downto 0);
Float149 : in STD_LOGIC_VECTOR (31 downto 0);
Float150 : in STD_LOGIC_VECTOR (31 downto 0);
Somme_out : out STD_LOGIC_VECTOR (31 downto 0));
end W150_Adder;

Architecture Behavioral of W150_Adder is

signal RAM_Out001 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out002 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out003 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out004 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out005 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out006 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out007 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out008 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out009 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out010 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out011 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out012 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out013 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out014 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out015 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out016 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out017 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out018 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out019 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out020 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out021 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out022 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out023 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out024 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out025 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out026 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out027 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out028 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out029 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out030 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out031 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out032 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out033 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out034 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out035 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out036 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out037 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out038 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out039 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out040 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out041 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out042 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out043 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out044 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out045 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out046 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out047 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out048 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out049 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out050 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out051 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out052 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out053 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out054 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out055 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out056 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out057 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out058 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out059 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out060 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out061 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out062 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out063 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out064 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out065 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out066 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out067 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out068 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out069 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out070 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out071 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out072 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out073 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out074 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out075 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out076 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out077 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out078 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out079 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out080 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out081 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out082 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out083 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out084 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out085 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out086 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out087 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out088 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out089 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out090 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out091 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out092 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out093 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out094 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out095 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out096 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out097 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out098 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out099 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out100 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out101 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out102 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out103 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out104 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out105 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out106 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out107 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out108 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out109 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out110 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out111 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out112 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out113 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out114 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out115 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out116 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out117 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out118 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out119 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out120 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out121 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out122 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out123 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out124 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out125 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out126 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out127 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out128 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out129 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out130 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out131 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out132 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out133 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out134 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out135 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out136 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out137 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out138 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out139 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out140 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out141 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out142 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out143 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out144 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out145 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out146 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out147 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out148 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out149 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Out150 : STD_LOGIC_VECTOR (31 downto 0);
signal RAM_Bias   : STD_LOGIC_VECTOR (31 downto 0);

signal Res_Mul001 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul002 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul003 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul004 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul005 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul006 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul007 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul008 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul009 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul010 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul011 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul012 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul013 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul014 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul015 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul016 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul017 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul018 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul019 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul020 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul021 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul022 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul023 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul024 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul025 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul026 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul027 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul028 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul029 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul030 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul031 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul032 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul033 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul034 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul035 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul036 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul037 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul038 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul039 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul040 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul041 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul042 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul043 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul044 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul045 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul046 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul047 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul048 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul049 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul050 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul051 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul052 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul053 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul054 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul055 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul056 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul057 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul058 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul059 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul060 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul061 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul062 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul063 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul064 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul065 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul066 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul067 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul068 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul069 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul070 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul071 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul072 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul073 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul074 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul075 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul076 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul077 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul078 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul079 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul080 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul081 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul082 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul083 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul084 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul085 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul086 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul087 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul088 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul089 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul090 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul091 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul092 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul093 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul094 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul095 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul096 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul097 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul098 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul099 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul100 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul101 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul102 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul103 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul104 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul105 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul106 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul107 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul108 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul109 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul110 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul111 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul112 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul113 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul114 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul115 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul116 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul117 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul118 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul119 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul120 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul121 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul122 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul123 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul124 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul125 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul126 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul127 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul128 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul129 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul130 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul131 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul132 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul133 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul134 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul135 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul136 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul137 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul138 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul139 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul140 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul141 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul142 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul143 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul144 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul145 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul146 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul147 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul148 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul149 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Mul150 : STD_LOGIC_VECTOR (31 downto 0);

signal Res_Adder001 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder002 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder003 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder004 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder005 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder006 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder007 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder008 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder009 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder010 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder011 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder012 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder013 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder014 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder015 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder016 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder017 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder018 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder019 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder020 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder021 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder022 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder023 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder024 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder025 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder026 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder027 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder028 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder029 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder030 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder031 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder032 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder033 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder034 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder035 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder036 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder037 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder038 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder039 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder040 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder041 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder042 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder043 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder044 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder045 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder046 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder047 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder048 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder049 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder050 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder051 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder052 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder053 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder054 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder055 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder056 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder057 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder058 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder059 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder060 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder061 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder062 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder063 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder064 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder065 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder066 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder067 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder068 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder069 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder070 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder071 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder072 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder073 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder074 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder075 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder076 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder077 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder078 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder079 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder080 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder081 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder082 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder083 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder084 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder085 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder086 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder087 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder088 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder089 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder090 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder091 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder092 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder093 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder094 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder095 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder096 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder097 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder098 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder099 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder100 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder101 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder102 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder103 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder104 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder105 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder106 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder107 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder108 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder109 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder110 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder111 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder112 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder113 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder114 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder115 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder116 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder117 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder118 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder119 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder120 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder121 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder122 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder123 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder124 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder125 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder126 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder127 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder128 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder129 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder130 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder131 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder132 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder133 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder134 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder135 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder136 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder137 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder138 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder139 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder140 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder141 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder142 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder143 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder144 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder145 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder146 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder147 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder148 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder149 : STD_LOGIC_VECTOR (31 downto 0);
signal Res_Adder150 : STD_LOGIC_VECTOR (31 downto 0);

Component multiplier_organised is
Port ( x : in  STD_LOGIC_VECTOR (31 downto 0);
       y : in  STD_LOGIC_VECTOR (31 downto 0);
       z : out STD_LOGIC_VECTOR (31 downto 0));
end Component;

Component adder_single_precision is
    Port (  CLK, RST :      in  STD_LOGIC;
            Float1, Float2: in  STD_LOGIC_vector(31 downto 0);
            output :        out STD_LOGIC_vector(31 downto 0));
end Component;

begin

    Mul001 : multiplier_organised port map (Float001, RAM_Out001, Res_Mul001);
    Mul002 : multiplier_organised port map (Float002, RAM_Out002, Res_Mul002);
    Mul003 : multiplier_organised port map (Float003, RAM_Out003, Res_Mul003);
    Mul004 : multiplier_organised port map (Float004, RAM_Out004, Res_Mul004);
    Mul005 : multiplier_organised port map (Float005, RAM_Out005, Res_Mul005);
    Mul006 : multiplier_organised port map (Float006, RAM_Out006, Res_Mul006);
    Mul007 : multiplier_organised port map (Float007, RAM_Out007, Res_Mul007);
    Mul008 : multiplier_organised port map (Float008, RAM_Out008, Res_Mul008);
    Mul009 : multiplier_organised port map (Float009, RAM_Out009, Res_Mul009);
    Mul010 : multiplier_organised port map (Float010, RAM_Out010, Res_Mul010);
    Mul011 : multiplier_organised port map (Float011, RAM_Out011, Res_Mul011);
    Mul012 : multiplier_organised port map (Float012, RAM_Out012, Res_Mul012);
    Mul013 : multiplier_organised port map (Float013, RAM_Out013, Res_Mul013);
    Mul014 : multiplier_organised port map (Float014, RAM_Out014, Res_Mul014);
    Mul015 : multiplier_organised port map (Float015, RAM_Out015, Res_Mul015);
    Mul016 : multiplier_organised port map (Float016, RAM_Out016, Res_Mul016);
    Mul017 : multiplier_organised port map (Float017, RAM_Out017, Res_Mul017);
    Mul018 : multiplier_organised port map (Float018, RAM_Out018, Res_Mul018);
    Mul019 : multiplier_organised port map (Float019, RAM_Out019, Res_Mul019);
    Mul020 : multiplier_organised port map (Float020, RAM_Out020, Res_Mul020);
    Mul021 : multiplier_organised port map (Float021, RAM_Out021, Res_Mul021);
    Mul022 : multiplier_organised port map (Float022, RAM_Out022, Res_Mul022);
    Mul023 : multiplier_organised port map (Float023, RAM_Out023, Res_Mul023);
    Mul024 : multiplier_organised port map (Float024, RAM_Out024, Res_Mul024);
    Mul025 : multiplier_organised port map (Float025, RAM_Out025, Res_Mul025);
    Mul026 : multiplier_organised port map (Float026, RAM_Out026, Res_Mul026);
    Mul027 : multiplier_organised port map (Float027, RAM_Out027, Res_Mul027);
    Mul028 : multiplier_organised port map (Float028, RAM_Out028, Res_Mul028);
    Mul029 : multiplier_organised port map (Float029, RAM_Out029, Res_Mul029);
    Mul030 : multiplier_organised port map (Float030, RAM_Out030, Res_Mul030);
    Mul031 : multiplier_organised port map (Float031, RAM_Out031, Res_Mul031);
    Mul032 : multiplier_organised port map (Float032, RAM_Out032, Res_Mul032);
    Mul033 : multiplier_organised port map (Float033, RAM_Out033, Res_Mul033);
    Mul034 : multiplier_organised port map (Float034, RAM_Out034, Res_Mul034);
    Mul035 : multiplier_organised port map (Float035, RAM_Out035, Res_Mul035);
    Mul036 : multiplier_organised port map (Float036, RAM_Out036, Res_Mul036);
    Mul037 : multiplier_organised port map (Float037, RAM_Out037, Res_Mul037);
    Mul038 : multiplier_organised port map (Float038, RAM_Out038, Res_Mul038);
    Mul039 : multiplier_organised port map (Float039, RAM_Out039, Res_Mul039);
    Mul040 : multiplier_organised port map (Float040, RAM_Out040, Res_Mul040);
    Mul041 : multiplier_organised port map (Float041, RAM_Out041, Res_Mul041);
    Mul042 : multiplier_organised port map (Float042, RAM_Out042, Res_Mul042);
    Mul043 : multiplier_organised port map (Float043, RAM_Out043, Res_Mul043);
    Mul044 : multiplier_organised port map (Float044, RAM_Out044, Res_Mul044);
    Mul045 : multiplier_organised port map (Float045, RAM_Out045, Res_Mul045);
    Mul046 : multiplier_organised port map (Float046, RAM_Out046, Res_Mul046);
    Mul047 : multiplier_organised port map (Float047, RAM_Out047, Res_Mul047);
    Mul048 : multiplier_organised port map (Float048, RAM_Out048, Res_Mul048);
    Mul049 : multiplier_organised port map (Float049, RAM_Out049, Res_Mul049);
    Mul050 : multiplier_organised port map (Float050, RAM_Out050, Res_Mul050);
    Mul051 : multiplier_organised port map (Float051, RAM_Out051, Res_Mul051);
    Mul052 : multiplier_organised port map (Float052, RAM_Out052, Res_Mul052);
    Mul053 : multiplier_organised port map (Float053, RAM_Out053, Res_Mul053);
    Mul054 : multiplier_organised port map (Float054, RAM_Out054, Res_Mul054);
    Mul055 : multiplier_organised port map (Float055, RAM_Out055, Res_Mul055);
    Mul056 : multiplier_organised port map (Float056, RAM_Out056, Res_Mul056);
    Mul057 : multiplier_organised port map (Float057, RAM_Out057, Res_Mul057);
    Mul058 : multiplier_organised port map (Float058, RAM_Out058, Res_Mul058);
    Mul059 : multiplier_organised port map (Float059, RAM_Out059, Res_Mul059);
    Mul060 : multiplier_organised port map (Float060, RAM_Out060, Res_Mul060);
    Mul061 : multiplier_organised port map (Float061, RAM_Out061, Res_Mul061);
    Mul062 : multiplier_organised port map (Float062, RAM_Out062, Res_Mul062);
    Mul063 : multiplier_organised port map (Float063, RAM_Out063, Res_Mul063);
    Mul064 : multiplier_organised port map (Float064, RAM_Out064, Res_Mul064);
    Mul065 : multiplier_organised port map (Float065, RAM_Out065, Res_Mul065);
    Mul066 : multiplier_organised port map (Float066, RAM_Out066, Res_Mul066);
    Mul067 : multiplier_organised port map (Float067, RAM_Out067, Res_Mul067);
    Mul068 : multiplier_organised port map (Float068, RAM_Out068, Res_Mul068);
    Mul069 : multiplier_organised port map (Float069, RAM_Out069, Res_Mul069);
    Mul070 : multiplier_organised port map (Float070, RAM_Out070, Res_Mul070);
    Mul071 : multiplier_organised port map (Float071, RAM_Out071, Res_Mul071);
    Mul072 : multiplier_organised port map (Float072, RAM_Out072, Res_Mul072);
    Mul073 : multiplier_organised port map (Float073, RAM_Out073, Res_Mul073);
    Mul074 : multiplier_organised port map (Float074, RAM_Out074, Res_Mul074);
    Mul075 : multiplier_organised port map (Float075, RAM_Out075, Res_Mul075);
    Mul076 : multiplier_organised port map (Float076, RAM_Out076, Res_Mul076);
    Mul077 : multiplier_organised port map (Float077, RAM_Out077, Res_Mul077);
    Mul078 : multiplier_organised port map (Float078, RAM_Out078, Res_Mul078);
    Mul079 : multiplier_organised port map (Float079, RAM_Out079, Res_Mul079);
    Mul080 : multiplier_organised port map (Float080, RAM_Out080, Res_Mul080);
    Mul081 : multiplier_organised port map (Float081, RAM_Out081, Res_Mul081);
    Mul082 : multiplier_organised port map (Float082, RAM_Out082, Res_Mul082);
    Mul083 : multiplier_organised port map (Float083, RAM_Out083, Res_Mul083);
    Mul084 : multiplier_organised port map (Float084, RAM_Out084, Res_Mul084);
    Mul085 : multiplier_organised port map (Float085, RAM_Out085, Res_Mul085);
    Mul086 : multiplier_organised port map (Float086, RAM_Out086, Res_Mul086);
    Mul087 : multiplier_organised port map (Float087, RAM_Out087, Res_Mul087);
    Mul088 : multiplier_organised port map (Float088, RAM_Out088, Res_Mul088);
    Mul089 : multiplier_organised port map (Float089, RAM_Out089, Res_Mul089);
    Mul090 : multiplier_organised port map (Float090, RAM_Out090, Res_Mul090);
    Mul091 : multiplier_organised port map (Float091, RAM_Out091, Res_Mul091);
    Mul092 : multiplier_organised port map (Float092, RAM_Out092, Res_Mul092);
    Mul093 : multiplier_organised port map (Float093, RAM_Out093, Res_Mul093);
    Mul094 : multiplier_organised port map (Float094, RAM_Out094, Res_Mul094);
    Mul095 : multiplier_organised port map (Float095, RAM_Out095, Res_Mul095);
    Mul096 : multiplier_organised port map (Float096, RAM_Out096, Res_Mul096);
    Mul097 : multiplier_organised port map (Float097, RAM_Out097, Res_Mul097);
    Mul098 : multiplier_organised port map (Float098, RAM_Out098, Res_Mul098);
    Mul099 : multiplier_organised port map (Float099, RAM_Out099, Res_Mul099);
    Mul100 : multiplier_organised port map (Float100, RAM_Out100, Res_Mul100);
    Mul101 : multiplier_organised port map (Float101, RAM_Out101, Res_Mul101);
    Mul102 : multiplier_organised port map (Float102, RAM_Out102, Res_Mul102);
    Mul103 : multiplier_organised port map (Float103, RAM_Out103, Res_Mul103);
    Mul104 : multiplier_organised port map (Float104, RAM_Out104, Res_Mul104);
    Mul105 : multiplier_organised port map (Float105, RAM_Out105, Res_Mul105);
    Mul106 : multiplier_organised port map (Float106, RAM_Out106, Res_Mul106);
    Mul107 : multiplier_organised port map (Float107, RAM_Out107, Res_Mul107);
    Mul108 : multiplier_organised port map (Float108, RAM_Out108, Res_Mul108);
    Mul109 : multiplier_organised port map (Float109, RAM_Out109, Res_Mul109);
    Mul110 : multiplier_organised port map (Float110, RAM_Out110, Res_Mul110);
    Mul111 : multiplier_organised port map (Float111, RAM_Out111, Res_Mul111);
    Mul112 : multiplier_organised port map (Float112, RAM_Out112, Res_Mul112);
    Mul113 : multiplier_organised port map (Float113, RAM_Out113, Res_Mul113);
    Mul114 : multiplier_organised port map (Float114, RAM_Out114, Res_Mul114);
    Mul115 : multiplier_organised port map (Float115, RAM_Out115, Res_Mul115);
    Mul116 : multiplier_organised port map (Float116, RAM_Out116, Res_Mul116);
    Mul117 : multiplier_organised port map (Float117, RAM_Out117, Res_Mul117);
    Mul118 : multiplier_organised port map (Float118, RAM_Out118, Res_Mul118);
    Mul119 : multiplier_organised port map (Float119, RAM_Out119, Res_Mul119);
    Mul120 : multiplier_organised port map (Float120, RAM_Out120, Res_Mul120);
    Mul121 : multiplier_organised port map (Float121, RAM_Out121, Res_Mul121);
    Mul122 : multiplier_organised port map (Float122, RAM_Out122, Res_Mul122);
    Mul123 : multiplier_organised port map (Float123, RAM_Out123, Res_Mul123);
    Mul124 : multiplier_organised port map (Float124, RAM_Out124, Res_Mul124);
    Mul125 : multiplier_organised port map (Float125, RAM_Out125, Res_Mul125);
    Mul126 : multiplier_organised port map (Float126, RAM_Out126, Res_Mul126);
    Mul127 : multiplier_organised port map (Float127, RAM_Out127, Res_Mul127);
    Mul128 : multiplier_organised port map (Float128, RAM_Out128, Res_Mul128);
    Mul129 : multiplier_organised port map (Float129, RAM_Out129, Res_Mul129);
    Mul130 : multiplier_organised port map (Float130, RAM_Out130, Res_Mul130);
    Mul131 : multiplier_organised port map (Float131, RAM_Out131, Res_Mul131);
    Mul132 : multiplier_organised port map (Float132, RAM_Out132, Res_Mul132);
    Mul133 : multiplier_organised port map (Float133, RAM_Out133, Res_Mul133);
    Mul134 : multiplier_organised port map (Float134, RAM_Out134, Res_Mul134);
    Mul135 : multiplier_organised port map (Float135, RAM_Out135, Res_Mul135);
    Mul136 : multiplier_organised port map (Float136, RAM_Out136, Res_Mul136);
    Mul137 : multiplier_organised port map (Float137, RAM_Out137, Res_Mul137);
    Mul138 : multiplier_organised port map (Float138, RAM_Out138, Res_Mul138);
    Mul139 : multiplier_organised port map (Float139, RAM_Out139, Res_Mul139);
    Mul140 : multiplier_organised port map (Float140, RAM_Out140, Res_Mul140);
    Mul141 : multiplier_organised port map (Float141, RAM_Out141, Res_Mul141);
    Mul142 : multiplier_organised port map (Float142, RAM_Out142, Res_Mul142);
    Mul143 : multiplier_organised port map (Float143, RAM_Out143, Res_Mul143);
    Mul144 : multiplier_organised port map (Float144, RAM_Out144, Res_Mul144);
    Mul145 : multiplier_organised port map (Float145, RAM_Out145, Res_Mul145);
    Mul146 : multiplier_organised port map (Float146, RAM_Out146, Res_Mul146);
    Mul147 : multiplier_organised port map (Float147, RAM_Out147, Res_Mul147);
    Mul148 : multiplier_organised port map (Float148, RAM_Out148, Res_Mul148);
    Mul149 : multiplier_organised port map (Float149, RAM_Out149, Res_Mul149);
    Mul150 : multiplier_organised port map (Float150, RAM_Out150, Res_Mul150);

    Adder001 : adder_single_precision port map (CLK, RST, Res_Mul001, Res_Mul002, Res_Adder001);
    Adder002 : adder_single_precision port map (CLK, RST, Res_Mul003, Res_Mul004, Res_Adder002);
    Adder003 : adder_single_precision port map (CLK, RST, Res_Mul005, Res_Mul006, Res_Adder003);
    Adder004 : adder_single_precision port map (CLK, RST, Res_Mul007, Res_Mul008, Res_Adder004);
    Adder005 : adder_single_precision port map (CLK, RST, Res_Mul009, Res_Mul150, Res_Adder005);
    Adder006 : adder_single_precision port map (CLK, RST, Res_Mul011, Res_Mul012, Res_Adder006);
    Adder007 : adder_single_precision port map (CLK, RST, Res_Mul013, Res_Mul014, Res_Adder007);
    Adder008 : adder_single_precision port map (CLK, RST, Res_Mul015, Res_Mul016, Res_Adder008);
    Adder009 : adder_single_precision port map (CLK, RST, Res_Mul017, Res_Mul018, Res_Adder009);
    Adder010 : adder_single_precision port map (CLK, RST, Res_Mul019, Res_Mul010, Res_Adder010);
    Adder011 : adder_single_precision port map (CLK, RST, Res_Mul021, Res_Mul022, Res_Adder011);
    Adder012 : adder_single_precision port map (CLK, RST, Res_Mul023, Res_Mul024, Res_Adder012);
    Adder013 : adder_single_precision port map (CLK, RST, Res_Mul025, Res_Mul026, Res_Adder013);
    Adder014 : adder_single_precision port map (CLK, RST, Res_Mul027, Res_Mul028, Res_Adder014);
    Adder015 : adder_single_precision port map (CLK, RST, Res_Mul029, Res_Mul020, Res_Adder015);
    Adder016 : adder_single_precision port map (CLK, RST, Res_Mul031, Res_Mul032, Res_Adder016);
    Adder017 : adder_single_precision port map (CLK, RST, Res_Mul033, Res_Mul034, Res_Adder017);
    Adder018 : adder_single_precision port map (CLK, RST, Res_Mul035, Res_Mul036, Res_Adder018);
    Adder019 : adder_single_precision port map (CLK, RST, Res_Mul037, Res_Mul038, Res_Adder019);
    Adder020 : adder_single_precision port map (CLK, RST, Res_Mul039, Res_Mul030, Res_Adder020);
    Adder021 : adder_single_precision port map (CLK, RST, Res_Mul041, Res_Mul042, Res_Adder021);
    Adder022 : adder_single_precision port map (CLK, RST, Res_Mul043, Res_Mul044, Res_Adder022);
    Adder023 : adder_single_precision port map (CLK, RST, Res_Mul045, Res_Mul046, Res_Adder023);
    Adder024 : adder_single_precision port map (CLK, RST, Res_Mul047, Res_Mul048, Res_Adder024);
    Adder025 : adder_single_precision port map (CLK, RST, Res_Mul049, Res_Mul040, Res_Adder025);
    Adder026 : adder_single_precision port map (CLK, RST, Res_Mul051, Res_Mul052, Res_Adder026);
    Adder027 : adder_single_precision port map (CLK, RST, Res_Mul053, Res_Mul054, Res_Adder027);
    Adder028 : adder_single_precision port map (CLK, RST, Res_Mul055, Res_Mul056, Res_Adder028);
    Adder029 : adder_single_precision port map (CLK, RST, Res_Mul057, Res_Mul058, Res_Adder029);
    Adder030 : adder_single_precision port map (CLK, RST, Res_Mul059, Res_Mul050, Res_Adder030);
    Adder031 : adder_single_precision port map (CLK, RST, Res_Mul061, Res_Mul062, Res_Adder031);
    Adder032 : adder_single_precision port map (CLK, RST, Res_Mul063, Res_Mul064, Res_Adder032);
    Adder033 : adder_single_precision port map (CLK, RST, Res_Mul065, Res_Mul066, Res_Adder033);
    Adder034 : adder_single_precision port map (CLK, RST, Res_Mul067, Res_Mul068, Res_Adder034);
    Adder035 : adder_single_precision port map (CLK, RST, Res_Mul069, Res_Mul060, Res_Adder035);
    Adder036 : adder_single_precision port map (CLK, RST, Res_Mul071, Res_Mul072, Res_Adder036);
    Adder037 : adder_single_precision port map (CLK, RST, Res_Mul073, Res_Mul074, Res_Adder037);
    Adder038 : adder_single_precision port map (CLK, RST, Res_Mul075, Res_Mul076, Res_Adder038);
    Adder039 : adder_single_precision port map (CLK, RST, Res_Mul077, Res_Mul078, Res_Adder039);
    Adder040 : adder_single_precision port map (CLK, RST, Res_Mul079, Res_Mul070, Res_Adder040);
    Adder041 : adder_single_precision port map (CLK, RST, Res_Mul081, Res_Mul082, Res_Adder041);
    Adder042 : adder_single_precision port map (CLK, RST, Res_Mul083, Res_Mul084, Res_Adder042);
    Adder043 : adder_single_precision port map (CLK, RST, Res_Mul085, Res_Mul086, Res_Adder043);
    Adder044 : adder_single_precision port map (CLK, RST, Res_Mul087, Res_Mul088, Res_Adder044);
    Adder045 : adder_single_precision port map (CLK, RST, Res_Mul089, Res_Mul080, Res_Adder045);
    Adder046 : adder_single_precision port map (CLK, RST, Res_Mul091, Res_Mul092, Res_Adder046);
    Adder047 : adder_single_precision port map (CLK, RST, Res_Mul093, Res_Mul094, Res_Adder047);
    Adder048 : adder_single_precision port map (CLK, RST, Res_Mul095, Res_Mul096, Res_Adder048);
    Adder049 : adder_single_precision port map (CLK, RST, Res_Mul097, Res_Mul098, Res_Adder049);
    Adder050 : adder_single_precision port map (CLK, RST, Res_Mul099, Res_Mul090, Res_Adder050);
    Adder051 : adder_single_precision port map (CLK, RST, Res_Mul101, Res_Mul102, Res_Adder051);
    Adder052 : adder_single_precision port map (CLK, RST, Res_Mul103, Res_Mul104, Res_Adder052);
    Adder053 : adder_single_precision port map (CLK, RST, Res_Mul105, Res_Mul106, Res_Adder053);
    Adder054 : adder_single_precision port map (CLK, RST, Res_Mul107, Res_Mul108, Res_Adder054);
    Adder055 : adder_single_precision port map (CLK, RST, Res_Mul109, Res_Mul100, Res_Adder055);
    Adder056 : adder_single_precision port map (CLK, RST, Res_Mul111, Res_Mul112, Res_Adder056);
    Adder057 : adder_single_precision port map (CLK, RST, Res_Mul113, Res_Mul114, Res_Adder057);
    Adder058 : adder_single_precision port map (CLK, RST, Res_Mul115, Res_Mul116, Res_Adder058);
    Adder059 : adder_single_precision port map (CLK, RST, Res_Mul117, Res_Mul118, Res_Adder059);
    Adder060 : adder_single_precision port map (CLK, RST, Res_Mul119, Res_Mul110, Res_Adder060);
    Adder061 : adder_single_precision port map (CLK, RST, Res_Mul121, Res_Mul122, Res_Adder061);
    Adder062 : adder_single_precision port map (CLK, RST, Res_Mul123, Res_Mul124, Res_Adder062);
    Adder063 : adder_single_precision port map (CLK, RST, Res_Mul125, Res_Mul126, Res_Adder063);
    Adder064 : adder_single_precision port map (CLK, RST, Res_Mul127, Res_Mul128, Res_Adder064);
    Adder065 : adder_single_precision port map (CLK, RST, Res_Mul129, Res_Mul120, Res_Adder065);
    Adder066 : adder_single_precision port map (CLK, RST, Res_Mul131, Res_Mul132, Res_Adder066);
    Adder067 : adder_single_precision port map (CLK, RST, Res_Mul133, Res_Mul134, Res_Adder067);
    Adder068 : adder_single_precision port map (CLK, RST, Res_Mul135, Res_Mul136, Res_Adder068);
    Adder069 : adder_single_precision port map (CLK, RST, Res_Mul137, Res_Mul138, Res_Adder069);
    Adder070 : adder_single_precision port map (CLK, RST, Res_Mul139, Res_Mul130, Res_Adder070);
    Adder071 : adder_single_precision port map (CLK, RST, Res_Mul141, Res_Mul142, Res_Adder071);
    Adder072 : adder_single_precision port map (CLK, RST, Res_Mul143, Res_Mul144, Res_Adder072);
    Adder073 : adder_single_precision port map (CLK, RST, Res_Mul145, Res_Mul146, Res_Adder073);
    Adder074 : adder_single_precision port map (CLK, RST, Res_Mul147, Res_Mul148, Res_Adder074);
    Adder075 : adder_single_precision port map (CLK, RST, Res_Mul149, Res_Mul140, Res_Adder075);
    Adder076 : adder_single_precision port map (CLK, RST, Res_Adder001, Res_Adder002, Res_Adder076);
    Adder077 : adder_single_precision port map (CLK, RST, Res_Adder003, Res_Adder004, Res_Adder077);
    Adder078 : adder_single_precision port map (CLK, RST, Res_Adder005, Res_Adder006, Res_Adder078);
    Adder079 : adder_single_precision port map (CLK, RST, Res_Adder007, Res_Adder008, Res_Adder079);
    Adder080 : adder_single_precision port map (CLK, RST, Res_Adder009, Res_Adder010, Res_Adder080);
    Adder081 : adder_single_precision port map (CLK, RST, Res_Adder011, Res_Adder012, Res_Adder081);
    Adder082 : adder_single_precision port map (CLK, RST, Res_Adder013, Res_Adder014, Res_Adder082);
    Adder083 : adder_single_precision port map (CLK, RST, Res_Adder015, Res_Adder016, Res_Adder083);
    Adder084 : adder_single_precision port map (CLK, RST, Res_Adder017, Res_Adder018, Res_Adder084);
    Adder085 : adder_single_precision port map (CLK, RST, Res_Adder019, Res_Adder020, Res_Adder085);
    Adder086 : adder_single_precision port map (CLK, RST, Res_Adder021, Res_Adder022, Res_Adder086);
    Adder087 : adder_single_precision port map (CLK, RST, Res_Adder023, Res_Adder024, Res_Adder087);
    Adder088 : adder_single_precision port map (CLK, RST, Res_Adder025, Res_Adder026, Res_Adder088);
    Adder089 : adder_single_precision port map (CLK, RST, Res_Adder027, Res_Adder028, Res_Adder089);
    Adder090 : adder_single_precision port map (CLK, RST, Res_Adder029, Res_Adder030, Res_Adder090);
    Adder091 : adder_single_precision port map (CLK, RST, Res_Adder031, Res_Adder032, Res_Adder091);
    Adder092 : adder_single_precision port map (CLK, RST, Res_Adder033, Res_Adder034, Res_Adder092);
    Adder093 : adder_single_precision port map (CLK, RST, Res_Adder035, Res_Adder036, Res_Adder093);
    Adder094 : adder_single_precision port map (CLK, RST, Res_Adder037, Res_Adder038, Res_Adder094);
    Adder095 : adder_single_precision port map (CLK, RST, Res_Adder039, Res_Adder040, Res_Adder095);
    Adder096 : adder_single_precision port map (CLK, RST, Res_Adder041, Res_Adder042, Res_Adder096);
    Adder097 : adder_single_precision port map (CLK, RST, Res_Adder043, Res_Adder044, Res_Adder097);
    Adder098 : adder_single_precision port map (CLK, RST, Res_Adder045, Res_Adder046, Res_Adder098);
    Adder099 : adder_single_precision port map (CLK, RST, Res_Adder047, Res_Adder048, Res_Adder099);
    Adder100 : adder_single_precision port map (CLK, RST, Res_Adder049, Res_Adder050, Res_Adder100);
    Adder101 : adder_single_precision port map (CLK, RST, Res_Adder051, Res_Adder052, Res_Adder101);
    Adder102 : adder_single_precision port map (CLK, RST, Res_Adder053, Res_Adder054, Res_Adder102);
    Adder103 : adder_single_precision port map (CLK, RST, Res_Adder055, Res_Adder056, Res_Adder103);
    Adder104 : adder_single_precision port map (CLK, RST, Res_Adder057, Res_Adder058, Res_Adder104);
    Adder105 : adder_single_precision port map (CLK, RST, Res_Adder059, Res_Adder060, Res_Adder105);
    Adder106 : adder_single_precision port map (CLK, RST, Res_Adder061, Res_Adder062, Res_Adder106);
    Adder107 : adder_single_precision port map (CLK, RST, Res_Adder063, Res_Adder064, Res_Adder107);
    Adder108 : adder_single_precision port map (CLK, RST, Res_Adder065, Res_Adder066, Res_Adder108);
    Adder109 : adder_single_precision port map (CLK, RST, Res_Adder067, Res_Adder068, Res_Adder109);
    Adder110 : adder_single_precision port map (CLK, RST, Res_Adder069, Res_Adder070, Res_Adder110);
    Adder111 : adder_single_precision port map (CLK, RST, Res_Adder071, Res_Adder072, Res_Adder111);
    Adder112 : adder_single_precision port map (CLK, RST, Res_Adder073, Res_Adder074, Res_Adder112);
    Adder113 : adder_single_precision port map (CLK, RST, Res_Adder075, Res_Adder076, Res_Adder113);
    Adder114 : adder_single_precision port map (CLK, RST, Res_Adder077, Res_Adder078, Res_Adder114);
    Adder115 : adder_single_precision port map (CLK, RST, Res_Adder079, Res_Adder080, Res_Adder115);
    Adder116 : adder_single_precision port map (CLK, RST, Res_Adder081, Res_Adder082, Res_Adder116);
    Adder117 : adder_single_precision port map (CLK, RST, Res_Adder083, Res_Adder084, Res_Adder117);
    Adder118 : adder_single_precision port map (CLK, RST, Res_Adder085, Res_Adder086, Res_Adder118);
    Adder119 : adder_single_precision port map (CLK, RST, Res_Adder087, Res_Adder088, Res_Adder119);
    Adder120 : adder_single_precision port map (CLK, RST, Res_Adder089, Res_Adder090, Res_Adder120);
    Adder121 : adder_single_precision port map (CLK, RST, Res_Adder091, Res_Adder092, Res_Adder121);
    Adder122 : adder_single_precision port map (CLK, RST, Res_Adder093, Res_Adder094, Res_Adder122);
    Adder123 : adder_single_precision port map (CLK, RST, Res_Adder095, Res_Adder096, Res_Adder123);
    Adder124 : adder_single_precision port map (CLK, RST, Res_Adder097, Res_Adder098, Res_Adder124);
    Adder125 : adder_single_precision port map (CLK, RST, Res_Adder099, Res_Adder100, Res_Adder125);
    Adder126 : adder_single_precision port map (CLK, RST, Res_Adder101, Res_Adder102, Res_Adder126);
    Adder127 : adder_single_precision port map (CLK, RST, Res_Adder103, Res_Adder104, Res_Adder127);
    Adder128 : adder_single_precision port map (CLK, RST, Res_Adder105, Res_Adder106, Res_Adder128);
    Adder129 : adder_single_precision port map (CLK, RST, Res_Adder107, Res_Adder108, Res_Adder129);
    Adder130 : adder_single_precision port map (CLK, RST, Res_Adder109, Res_Adder110, Res_Adder130);
    Adder131 : adder_single_precision port map (CLK, RST, Res_Adder111, Res_Adder112, Res_Adder131);
    Adder132 : adder_single_precision port map (CLK, RST, Res_Adder113, Res_Adder114, Res_Adder132);
    Adder133 : adder_single_precision port map (CLK, RST, Res_Adder115, Res_Adder116, Res_Adder133);
    Adder134 : adder_single_precision port map (CLK, RST, Res_Adder117, Res_Adder118, Res_Adder134);
    Adder135 : adder_single_precision port map (CLK, RST, Res_Adder119, Res_Adder120, Res_Adder135);
    Adder136 : adder_single_precision port map (CLK, RST, Res_Adder121, Res_Adder122, Res_Adder136);
    Adder137 : adder_single_precision port map (CLK, RST, Res_Adder123, Res_Adder124, Res_Adder137);
    Adder138 : adder_single_precision port map (CLK, RST, Res_Adder125, Res_Adder126, Res_Adder138);
    Adder139 : adder_single_precision port map (CLK, RST, Res_Adder127, Res_Adder128, Res_Adder139);
    Adder140 : adder_single_precision port map (CLK, RST, Res_Adder129, Res_Adder130, Res_Adder140);
    Adder141 : adder_single_precision port map (CLK, RST, Res_Adder131, Res_Adder132, Res_Adder141);
    Adder142 : adder_single_precision port map (CLK, RST, Res_Adder133, Res_Adder134, Res_Adder142);
    Adder143 : adder_single_precision port map (CLK, RST, Res_Adder135, Res_Adder136, Res_Adder143);
    Adder144 : adder_single_precision port map (CLK, RST, Res_Adder137, Res_Adder138, Res_Adder144);
    Adder145 : adder_single_precision port map (CLK, RST, Res_Adder139, Res_Adder140, Res_Adder145);
    Adder146 : adder_single_precision port map (CLK, RST, Res_Adder141, Res_Adder142, Res_Adder146);
    Adder147 : adder_single_precision port map (CLK, RST, Res_Adder143, Res_Adder144, Res_Adder147);
    Adder148 : adder_single_precision port map (CLK, RST, Res_Adder145, Res_Adder146, Res_Adder148);
    Adder149 : adder_single_precision port map (CLK, RST, Res_Adder147, Res_Adder148, Res_Adder149);
    Adder150 : adder_single_precision port map (CLK, RST, Res_Adder149, RAM_Bias, Res_Adder150);

    P1 : process(CLK, RST)
    begin
        if (WE = '1') then
            RAM_Bias   <= Bias;
            RAM_Out001 <= Float001;
            RAM_Out002 <= Float002;
            RAM_Out003 <= Float003;
            RAM_Out004 <= Float004;
            RAM_Out005 <= Float005;
            RAM_Out006 <= Float006;
            RAM_Out007 <= Float007;
            RAM_Out008 <= Float008;
            RAM_Out009 <= Float009;
            RAM_Out010 <= Float010;
            RAM_Out011 <= Float011;
            RAM_Out012 <= Float012;
            RAM_Out013 <= Float013;
            RAM_Out014 <= Float014;
            RAM_Out015 <= Float015;
            RAM_Out016 <= Float016;
            RAM_Out017 <= Float017;
            RAM_Out018 <= Float018;
            RAM_Out019 <= Float019;
            RAM_Out020 <= Float020;
            RAM_Out021 <= Float021;
            RAM_Out022 <= Float022;
            RAM_Out023 <= Float023;
            RAM_Out024 <= Float024;
            RAM_Out025 <= Float025;
            RAM_Out026 <= Float026;
            RAM_Out027 <= Float027;
            RAM_Out028 <= Float028;
            RAM_Out029 <= Float029;
            RAM_Out030 <= Float030;
            RAM_Out031 <= Float031;
            RAM_Out032 <= Float032;
            RAM_Out033 <= Float033;
            RAM_Out034 <= Float034;
            RAM_Out035 <= Float035;
            RAM_Out036 <= Float036;
            RAM_Out037 <= Float037;
            RAM_Out038 <= Float038;
            RAM_Out039 <= Float039;
            RAM_Out040 <= Float040;
            RAM_Out041 <= Float041;
            RAM_Out042 <= Float042;
            RAM_Out043 <= Float043;
            RAM_Out044 <= Float044;
            RAM_Out045 <= Float045;
            RAM_Out046 <= Float046;
            RAM_Out047 <= Float047;
            RAM_Out048 <= Float048;
            RAM_Out049 <= Float049;
            RAM_Out050 <= Float050;
            RAM_Out051 <= Float051;
            RAM_Out052 <= Float052;
            RAM_Out053 <= Float053;
            RAM_Out054 <= Float054;
            RAM_Out055 <= Float055;
            RAM_Out056 <= Float056;
            RAM_Out057 <= Float057;
            RAM_Out058 <= Float058;
            RAM_Out059 <= Float059;
            RAM_Out060 <= Float060;
            RAM_Out061 <= Float061;
            RAM_Out062 <= Float062;
            RAM_Out063 <= Float063;
            RAM_Out064 <= Float064;
            RAM_Out065 <= Float065;
            RAM_Out066 <= Float066;
            RAM_Out067 <= Float067;
            RAM_Out068 <= Float068;
            RAM_Out069 <= Float069;
            RAM_Out070 <= Float070;
            RAM_Out071 <= Float071;
            RAM_Out072 <= Float072;
            RAM_Out073 <= Float073;
            RAM_Out074 <= Float074;
            RAM_Out075 <= Float075;
            RAM_Out076 <= Float076;
            RAM_Out077 <= Float077;
            RAM_Out078 <= Float078;
            RAM_Out079 <= Float079;
            RAM_Out080 <= Float080;
            RAM_Out081 <= Float081;
            RAM_Out082 <= Float082;
            RAM_Out083 <= Float083;
            RAM_Out084 <= Float084;
            RAM_Out085 <= Float085;
            RAM_Out086 <= Float086;
            RAM_Out087 <= Float087;
            RAM_Out088 <= Float088;
            RAM_Out089 <= Float089;
            RAM_Out090 <= Float090;
            RAM_Out091 <= Float091;
            RAM_Out092 <= Float092;
            RAM_Out093 <= Float093;
            RAM_Out094 <= Float094;
            RAM_Out095 <= Float095;
            RAM_Out096 <= Float096;
            RAM_Out097 <= Float097;
            RAM_Out098 <= Float098;
            RAM_Out099 <= Float099;
            RAM_Out100 <= Float100;
            RAM_Out101 <= Float101;
            RAM_Out102 <= Float102;
            RAM_Out103 <= Float103;
            RAM_Out104 <= Float104;
            RAM_Out105 <= Float105;
            RAM_Out106 <= Float106;
            RAM_Out107 <= Float107;
            RAM_Out108 <= Float108;
            RAM_Out109 <= Float109;
            RAM_Out110 <= Float110;
            RAM_Out111 <= Float111;
            RAM_Out112 <= Float112;
            RAM_Out113 <= Float113;
            RAM_Out114 <= Float114;
            RAM_Out115 <= Float115;
            RAM_Out116 <= Float116;
            RAM_Out117 <= Float117;
            RAM_Out118 <= Float118;
            RAM_Out119 <= Float119;
            RAM_Out120 <= Float120;
            RAM_Out121 <= Float121;
            RAM_Out122 <= Float122;
            RAM_Out123 <= Float123;
            RAM_Out124 <= Float124;
            RAM_Out125 <= Float125;
            RAM_Out126 <= Float126;
            RAM_Out127 <= Float127;
            RAM_Out128 <= Float128;
            RAM_Out129 <= Float129;
            RAM_Out130 <= Float130;
            RAM_Out131 <= Float131;
            RAM_Out132 <= Float132;
            RAM_Out133 <= Float133;
            RAM_Out134 <= Float134;
            RAM_Out135 <= Float135;
            RAM_Out136 <= Float136;
            RAM_Out137 <= Float137;
            RAM_Out138 <= Float138;
            RAM_Out139 <= Float139;
            RAM_Out140 <= Float140;
            RAM_Out141 <= Float141;
            RAM_Out142 <= Float142;
            RAM_Out143 <= Float143;
            RAM_Out144 <= Float144;
            RAM_Out145 <= Float145;
            RAM_Out146 <= Float146;
            RAM_Out147 <= Float147;
            RAM_Out148 <= Float148;
            RAM_Out149 <= Float149;
            RAM_Out150 <= Float150;
        end if;
    end process P1;

    Somme_out <= Res_Adder150;

end Behavioral;
